`timescale 1ns / 1ps
`default_nettype none
`define OBJ_WIDTH 115
`define OBJ_COUNT 8
`define OBJ_ADDR_WIDTH 8
`define CLAMP(x, min, max) (x < min ? min : (x > max ? max : x))

module top_level
  (
    input wire          clk_100mhz,
    output logic [15:0] led,
    // camera bus
    input wire [7:0]    camera_d, // 8 parallel data wires
    output logic        cam_xclk, // XC driving camera
    input wire          cam_hsync, // camera hsync wire
    input wire          cam_vsync, // camera vsync wire
    input wire          cam_pclk, // camera pixel clock
    inout wire          i2c_scl, // i2c inout clock
    inout wire          i2c_sda, // i2c inout data
    input wire [15:0]   sw,
    input wire [3:0]    btn,
    output logic [2:0]  rgb0,
    output logic [2:0]  rgb1,
    // seven segment
    output logic [3:0]  ss0_an,//anode control for upper four digits of seven-seg display
    output logic [3:0]  ss1_an,//anode control for lower four digits of seven-seg display
    output logic [6:0]  ss0_c, //cathode controls for the segments of upper four digits
    output logic [6:0]  ss1_c, //cathod controls for the segments of lower four digits
    // hdmi port
    output logic [2:0]  hdmi_tx_p, //hdmi output signals (positives) (blue, green, red)
    output logic [2:0]  hdmi_tx_n, //hdmi output signals (negatives) (blue, green, red)
    output logic        hdmi_clk_p, hdmi_clk_n //differential hdmi clock
  );

  // shut up those RGBs
  assign rgb0 = 0;
  assign rgb1 = 0;

  // Clock and Reset Signals
  logic          sys_rst_camera;
  logic          sys_rst_pixel;

  logic          clk_camera;
  logic          clk_pixel;
  logic          clk_5x;
  logic          clk_xc;

  logic          clk_100_passthrough;

  // clocking wizards to generate the clock speeds we need for our different domains
  // clk_camera: 200MHz, fast enough to comfortably sample the cameera's PCLK (50MHz)
  cw_hdmi_clk_wiz wizard_hdmi
                  (.sysclk(clk_100_passthrough),
                   .clk_pixel(clk_pixel),
                   .clk_tmds(clk_5x),
                   .reset(0));

  cw_fast_clk_wiz wizard_migcam
                  (.clk_in1(clk_100mhz),
                   .clk_camera(clk_camera),
                   .clk_xc(clk_xc),
                   .clk_100(clk_100_passthrough),
                   .reset(0));

  // assign camera's xclk to pmod port: drive the operating clock of the camera!
  // this port also is specifically set to high drive by the XDC file.
  assign cam_xclk = sw[0] ? clk_xc : 1'b0;

  assign sys_rst_camera = btn[0]; //use for resetting camera side of logic
  assign sys_rst_pixel = btn[0]; //use for resetting hdmi/draw side of logic


  // video signal generator signals
  logic          hsync_hdmi;
  logic          vsync_hdmi;
  logic [10:0]  hcount_hdmi;
  logic [9:0]    vcount_hdmi;
  logic          active_draw_hdmi;
  logic          new_frame_hdmi;
  logic [5:0]    frame_count_hdmi;
  logic          nf_hdmi;

  // rgb output values
  logic [7:0]          red,green,blue;

  // ** Handling input from the camera **

  // synchronizers to prevent metastability
  logic [7:0]    camera_d_buf [1:0];
  logic          cam_hsync_buf [1:0];
  logic          cam_vsync_buf [1:0];
  logic          cam_pclk_buf [1:0];

  always_ff @(posedge clk_camera)
  begin
    camera_d_buf <= {camera_d, camera_d_buf[1]};
    cam_pclk_buf <= {cam_pclk, cam_pclk_buf[1]};
    cam_hsync_buf <= {cam_hsync, cam_hsync_buf[1]};
    cam_vsync_buf <= {cam_vsync, cam_vsync_buf[1]};
  end

  logic [10:0] camera_hcount;
  logic [9:0]  camera_vcount;
  logic [15:0] camera_pixel;
  logic        camera_valid;

  // your pixel_reconstruct module, from the exercise!
  // hook it up to buffered inputs.
  pixel_reconstruct pixel_constructor
    (.clk_in(clk_camera),
     .rst_in(sys_rst_camera),
     .camera_pclk_in(cam_pclk_buf[0]),
     .camera_hs_in(cam_hsync_buf[0]),
     .camera_vs_in(cam_vsync_buf[0]),
     .camera_data_in(camera_d_buf[0]),
     .pixel_valid_out(camera_valid),
     .pixel_hcount_out(camera_hcount),
     .pixel_vcount_out(camera_vcount),
     .pixel_data_out(camera_pixel));


  //two-port BRAM used to hold image from camera.
  //The camera is producing video at 720p and 30fps, but we can't store all of that
  //we're going to down-sample by a factor of 4 in both dimensions
  //so we have 320 by 180.  this is kinda a bummer, but we'll fix it
  //in future weeks by using off-chip DRAM.
  //even with the down-sample, because our camera is producing data at 30fps
  //and  our display is running at 720p at 60 fps, there's no hope to have the
  //production and consumption of information be synchronized in this system.
  //even if we could line it up once, the clocks of both systems will drift over time
  //so to avoid this sync issue, we use a conflict-resolution device...the frame buffer
  //instead we use a frame buffer as a go-between. The camera sends pixels in at
  //its own rate, and we pull them out for display at the 720p rate/requirement
  //this avoids the whole sync issue. It will however result in artifacts when you
  //introduce fast motion in front of the camera. These lines/tears in the image
  //are the result of unsynced frame-rewriting happening while displaying. It won't
  //matter for slow movement
  localparam FB_DEPTH = 320*180;
  localparam FB_SIZE = $clog2(FB_DEPTH);
  logic [FB_SIZE-1:0] addra; //used to specify address to write to in frame buffer

  logic valid_camera_mem; //used to enable writing pixel data to frame buffer
  logic [15:0] camera_mem; //used to pass pixel data into frame buffer


  //TO DO in camera part 1:
  always_ff @(posedge clk_camera)
  begin
    //create logic to handle wriiting of camera.
    //we want to down sample the data from the camera by a factor of four in both
    //the x and y dimensions! TO DO
    if (camera_valid)
    begin
      addra <= (camera_hcount) + ((camera_vcount) * 320);
      camera_mem <= camera_pixel;
      valid_camera_mem <= 1; // Enable memory write
    end
    else
    begin
      valid_camera_mem <= 0;
    end
  end

  //frame buffer from IP
  blk_mem_gen_0 frame_buffer (
                  .addra(addra), //pixels are stored using this math
                  .clka(clk_camera),
                  .wea(valid_camera_mem),
                  .dina(camera_mem),
                  .ena(1'b1),
                  .douta(), //never read from this side
                  .addrb(addrb),//transformed lookup pixel
                  .dinb(16'b0),
                  .clkb(clk_pixel),
                  .web(1'b0),
                  .enb(1'b1),
                  .doutb(frame_buff_raw)
                );
  logic [15:0] frame_buff_raw; //data out of frame buffer (565)
  logic [FB_SIZE-1:0] addrb; //used to lookup address in memory for reading from buffer
  logic good_addrb; //used to indicate within valid frame for scaling


  //TO DO in camera part 1:
  // Scale pixel coordinates from HDMI to the frame buffer to grab the right pixel
  //scaling logic!!! You need to complete!!! We want 1X, 2X, and 4X!
  always_ff @(posedge clk_pixel)
  begin
    //default: delete:
    // addrb <= (319-hcount_hdmi) + 320*vcount_hdmi;
    // good_addrb <= (hcount_hdmi<320)&&(vcount_hdmi<180);
    //use structure below to do scaling
    if (btn[1])
    begin //1X scaling from frame buffer
      addrb <= hcount_hdmi + vcount_hdmi * 320; //change me
      good_addrb <= (hcount_hdmi < 320) && (vcount_hdmi < 180); //change me
    end
    else if (!sw[0])
    begin //2X scaling from frame buffer
      addrb <= (hcount_hdmi >> 1) + (vcount_hdmi >> 1) * 320; //change me
      good_addrb <= (hcount_hdmi < 640) && (vcount_hdmi < 360); //change me
    end
    else
    begin //4X scaling from frame buffer
      addrb <= (hcount_hdmi >> 2) + (vcount_hdmi >> 2) * 320; // change me
      good_addrb <= (hcount_hdmi < 1280) && (vcount_hdmi < 720); //change me
    end
  end

  //split fame_buff into 3 8 bit color channels (5:6:5 adjusted accordingly)
  //remapped frame_buffer outputs with 8 bits for r, g, b
  logic [7:0] fb_red, fb_green, fb_blue;
  always_ff @(posedge clk_pixel)
  begin
    fb_red <= good_addrb?{frame_buff_raw[15:11],3'b0}:8'b0;
    fb_green <= good_addrb?{frame_buff_raw[10:5], 2'b0}:8'b0;
    fb_blue <= good_addrb?{frame_buff_raw[4:0],3'b0}:8'b0;
  end
  // Pixel Processing pre-HDMI output

  // RGB to YCrCb

  //output of rgb to ycrcb conversion (10 bits due to module):
  logic [9:0] y_full, cr_full, cb_full; //ycrcb conversion of full pixel
  //bottom 8 of y, cr, cb conversions:
  logic [7:0] y, cr, cb; //ycrcb conversion of full pixel
  //Convert RGB of full pixel to YCrCb
  //See lecture 07 for YCrCb discussion.
  //Module has a 3 cycle latency
  rgb_to_ycrcb rgbtoycrcb_m(
                 .clk_in(clk_pixel),
                 .r_in(fb_red),
                 .g_in(fb_green),
                 .b_in(fb_blue),
                 .y_out(y_full),
                 .cr_out(cr_full),
                 .cb_out(cb_full)
               );

  //channel select module (select which of six color channels to mask):
  // logic [2:0] channel_sel;
  logic [7:0] selected_channel; //selected channels
  //selected_channel could contain any of the six color channels depend on selection

  //threshold module (apply masking threshold):
  logic [7:0] lower_threshold;
  logic [7:0] upper_threshold;
  logic mask; //Whether or not thresholded pixel is 1 or 0

  //Center of Mass variables (tally all mask=1 pixels for a frame and calculate their center of mass)fb_red
  logic [10:0] x_com, x_com_calc; //long term x_com and output from module, resp
  logic [9:0] y_com, y_com_calc; //long term y_com and output from module, resp
  logic new_com; //used to know when to update x_com and y_com ...

  //channel select module (select which of six color channels to mask) FOR COM_2:
  // logic [2:0] channel_sel_2;
  logic [7:0] selected_channel_2; //selected channels
  //selected_channel could contain any of the six color channels depend on selection

  //threshold module (apply masking threshold) FOR COM_2:
  // logic [7:0] lower_threshold_2;
  // logic [7:0] upper_threshold_2;
  logic mask_2; //Whether or not thresholded pixel is 1 or 0

  //Center of Mass variables FOR COM_2 (tally all mask=1 pixels for a frame and calculate their center of mass)fb_red
  logic [10:0] x_com_2, x_com_calc_2; //long term x_com and output from module, resp
  logic [9:0] y_com_2, y_com_calc_2; //long term y_com and output from module, resp
  logic new_com_2; //used to know when to update x_com and y_com ...

  //take lower 8 of full outputs.
  // treat cr and cb as signed numbers, invert the MSB to get an unsigned equivalent ( [-128,128) maps to [0,256) )
  assign y = y_full[7:0];
  assign cr = {!cr_full[7],cr_full[6:0]};
  assign cb = {!cb_full[7],cb_full[6:0]};

  // PIPELINE LOGIC
  //vary the packed width based on signal
  //vary the unpacked width based on pipelining depth needed

  logic [7:0] fb_red_delayed_ps1;
  pipeline #(
             .WIDTH(8), .STAGES(3))
           fb_red_pipeline_ps1(
             .clk_pixel(clk_pixel),
             .signal(fb_red),
             //.stages(3),
             .delayed_signal(fb_red_delayed_ps1)
           );

  logic [7:0] fb_green_delayed_ps1;
  pipeline #(
             .WIDTH(8), .STAGES(3))
           fb_green_pipeline_ps1(
             .clk_pixel(clk_pixel),
             .signal(fb_green),
             //.stages(3),
             .delayed_signal(fb_green_delayed_ps1)
           );

  logic [7:0] fb_blue_delayed_ps1;
  pipeline #(
             .WIDTH(8), .STAGES(3))
           fb_blue_pipeline_ps1(
             .clk_pixel(clk_pixel),
             .signal(fb_blue),
             //.stages(3),
             .delayed_signal(fb_blue_delayed_ps1)
           );

  // assign channel_sel = 3'b101;

  // assign channel_sel_2 = 3'b110;
  // * 3'b000: green
  // * 3'b001: red
  // * 3'b010: blue
  // * 3'b011: not valid
  // * 3'b100: y (luminance)
  // * 3'b101: Cr (Chroma Red)
  // * 3'b110: Cb (Chroma Blue)
  // * 3'b111: not valid
  //Channel Select: Takes in the full RGB and YCrCb information and
  // chooses one of them to output as an 8 bit value
  // channel_select mcs(
  //    .sel_in(channel_sel),
  //    .r_in(fb_red_delayed_ps1),    //TODO: needs to use pipelined signal (PS1)
  //    .g_in(fb_green_delayed_ps1),  //TODO: needs to use pipelined signal (PS1)
  //    .b_in(fb_blue_delayed_ps1),   //TODO: needs to use pipelined signal (PS1)
  //    .y_in(y),
  //    .cr_in(cr),
  //    .cb_in(cb),
  //    .channel_out(selected_channel)
  // );

  // channel_select mcs_2(
  //    .sel_in(channel_sel_2),
  //    .r_in(fb_red_delayed_ps1),    //TODO: needs to use pipelined signal (PS1)
  //    .g_in(fb_green_delayed_ps1),  //TODO: needs to use pipelined signal (PS1)
  //    .b_in(fb_blue_delayed_ps1),   //TODO: needs to use pipelined signal (PS1)
  //    .y_in(y),
  //    .cr_in(cr),
  //    .cb_in(cb),
  //    .channel_out(selected_channel_2)
  // );

  assign selected_channel = cr;
  assign selected_channel_2 = cb;

  //threshold values used to determine what value  passes:
  assign lower_threshold = {4'b1010,4'b0};
  assign upper_threshold = {4'b1111,4'b0};
  //Thresholder: Takes in the full selected channedl and
  //based on upper and lower bounds provides a binary mask bit
  // * 1 if selected channel is within the bounds (inclusive)
  // * 0 if selected channel is not within the bounds
  threshold mt(
              .clk_in(clk_pixel),
              .rst_in(sys_rst_pixel),
              .pixel_in(selected_channel),
              .lower_bound_in(lower_threshold),
              .upper_bound_in(upper_threshold),
              .mask_out(mask) //single bit if pixel within mask.
            );

  threshold mt_2(
              .clk_in(clk_pixel),
              .rst_in(sys_rst_pixel),
              .pixel_in(selected_channel_2),
              .lower_bound_in(lower_threshold),
              .upper_bound_in(upper_threshold),
              .mask_out(mask_2) //single bit if pixel within mask.
            );

  // logic [26:0] nf_count;
  // evt_counter #(
  //       .MAX_COUNT(1280 * 720 >> 3)
  // ) count_nf(
  //       .clk_in(clk_pixel),
  //       .rst_in(sys_rst_pixel),
  //       .evt_in(nf_hdmi),
  //       .count_out(nf_count)
  //   );


  logic [6:0] cam_ss_c;
  logic [3:0] cam_ss0_an, cam_ss1_an;
  //modified version of seven segment display for showing
  // thresholds and selected channel
  // special customized version
  lab05_ssc mssc(.clk_in(clk_pixel),
                 .rst_in(sys_rst_pixel),
                 .lt_in(x_com),
                 .ut_in(x_com_2),
                 .channel_sel_in(3'b101),
                 .cat_out(cam_ss_c),
                 .an_out({cam_ss0_an, cam_ss1_an})
                );
  // assign ss0_c = ss_c; //control upper four digit's cathodes!
  // assign ss1_c = ss_c; //same as above but for lower four digits!
  assign ss0_c = simul_mode ? phys_ss_c : cam_ss_c;
  assign ss1_c = simul_mode ? phys_ss_c : cam_ss_c;
  assign ss0_an = simul_mode ? phys_ss0_an : cam_ss0_an;
  assign ss1_an = simul_mode ? phys_ss1_an : cam_ss1_an;

  logic [10:0] hcount_delayed_ps3;
  pipeline #(
             .WIDTH(11), .STAGES(8))
           hcount_pipeline_ps3(
             .clk_pixel(clk_pixel),
             .signal(hcount_hdmi),
             //.stages(8),
             .delayed_signal(hcount_delayed_ps3)
           );

  logic [9:0] vcount_delayed_ps3;
  pipeline #(
             .WIDTH(10), .STAGES(8))
           vcount_pipeline_ps3(
             .clk_pixel(clk_pixel),
             .signal(vcount_hdmi),
             //.stages(8),
             .delayed_signal(vcount_delayed_ps3)
           );

  logic nf_hdmi_delayed_ps3;
  pipeline #(
             .WIDTH(1), .STAGES(8))
           nf_hdmi_pipeline_ps3(
             .clk_pixel(clk_pixel),
             .signal(nf_hdmi),
             //.stages(8),
             .delayed_signal(nf_hdmi_delayed_ps3)
           );


  //Center of Mass Calculation: (you need to do)
  //using x_com_calc and y_com_calc values
  //Center of Mass:
  center_of_mass com_m(
                   .clk_in(clk_pixel),
                   .rst_in(sys_rst_pixel),
                   .x_in(hcount_delayed_ps3),  //TODO: needs to use pipelined signal! (PS3)
                   .y_in(vcount_delayed_ps3), //TODO: needs to use pipelined signal! (PS3)
                   .valid_in(mask), //aka threshold
                   .tabulate_in((nf_hdmi_delayed_ps3)),
                   .x_out(x_com_calc),
                   .y_out(y_com_calc),
                   .valid_out(new_com)
                 );

  center_of_mass com_m_2(
                   .clk_in(clk_pixel),
                   .rst_in(sys_rst_pixel),
                   .x_in(hcount_delayed_ps3),  //TODO: needs to use pipelined signal! (PS3)
                   .y_in(vcount_delayed_ps3), //TODO: needs to use pipelined signal! (PS3)
                   .valid_in(mask_2), //aka threshold
                   .tabulate_in((nf_hdmi_delayed_ps3)),
                   .x_out(x_com_calc_2),
                   .y_out(y_com_calc_2),
                   .valid_out(new_com_2)
                 );
  //grab logic for above
  //update center of mass x_com, y_com based on new_com signal
  always_ff @(posedge clk_pixel)
  begin
    if (sys_rst_pixel)
    begin
      x_com <= 0;
      y_com <= 0;
    end
    else if(new_com)
    begin
      x_com <= x_com_calc;
      y_com <= y_com_calc;
    end
    if (sys_rst_pixel)
    begin
      x_com_2 <= 0;
      y_com_2 <= 0;
    end
    else if(new_com_2)
    begin
      x_com_2 <= x_com_calc_2;
      y_com_2 <= y_com_calc_2;
    end
  end

  //rectangle output:
  logic in_rect;
  logic [83:0] rect_coord;
  logic rect_valid_out;

  //circle output:
  logic in_circle;
  logic [83:0] circle_coord;
  logic circle_valid_out;

  //line output:
  logic in_line;
  logic [83:0] line_coord;
  logic line_valid_out;

  logic [10:0] hcount_delayed_ps1;
  pipeline #(
             .WIDTH(11), .STAGES(3))
           hcount_pipeline_ps1(
             .clk_pixel(clk_pixel),
             .signal(hcount_hdmi),
             //.stages(3),
             .delayed_signal(hcount_delayed_ps1)
           );

  logic [9:0] vcount_delayed_ps1;
  pipeline #(
             .WIDTH(10), .STAGES(3))
           vcount_pipeline_ps1(
             .clk_pixel(clk_pixel),
             .signal(vcount_hdmi),
             //.stages(3),
             .delayed_signal(vcount_delayed_ps1)
           );

  draw_rectangle #(
                   .WIDTH(256),
                   .HEIGHT(256),
                   .COLOR(24'hFF_FF_FF))
                 rectangle (
                   .clk_in(clk_pixel),
                   .rst_in(sys_rst_pixel),
                   .valid_in(1),
                   .hcount_in(hcount_delayed_ps1),
                   .vcount_in(vcount_delayed_ps1),
                   .x_in_1(x_com),
                   .y_in_1(y_com),
                   .x_in_2(x_com_2),
                   .y_in_2(y_com_2),
                   .rect_coord(rect_coord),
                   .in_rect(in_rect),
                   .valid_out(rect_valid_out));


  draw_circle #(
                .WIDTH(256),
                .HEIGHT(256),
                .COLOR(24'hFF_FF_FF))
              circle (
                .clk_in(clk_pixel),
                .rst_in(sys_rst_pixel),
                .valid_in(1),
                .hcount_in(hcount_delayed_ps1),
                .vcount_in(vcount_delayed_ps1),
                .x_in_1(x_com),
                .y_in_1(y_com),
                .x_in_2(x_com_2),
                .y_in_2(y_com_2),
                .circle_coord(circle_coord),
                .in_circle(in_circle),
                .valid_out(circle_valid_out));

  draw_line #(
              .WIDTH(256),
              .HEIGHT(256),
              .COLOR(24'hFF_FF_FF))
            line (
              .clk_in(clk_pixel),
              .rst_in(sys_rst_pixel),
              .valid_in(1),
              .hcount_in(hcount_delayed_ps1),
              .vcount_in(vcount_delayed_ps1),
              .x_in_1(x_com),
              .y_in_1(y_com),
              .x_in_2(x_com_2),
              .y_in_2(y_com_2),
              .line_coord(line_coord),
              .in_line(in_line),
              .valid_out(line_valid_out));

  logic simul_mode;
  assign simul_mode = sw[15];


  // object storage RAM definition
  //  read from render and physics engine
  //  write from draw and physics engine

  logic write_valid_in;
  logic [`OBJ_ADDR_WIDTH-1:0] write_addr_in;
  logic [`OBJ_WIDTH-1:0] write_object_in;
  logic write_valid_out;

  logic read_valid_in;
  logic [`OBJ_ADDR_WIDTH-1:0] read_addrs_in [3:0];
  logic [`OBJ_WIDTH-1:0] read_objects_out [3:0];
  logic read_valid_out;

  object_storage storage(
                   .clk_in(clk_pixel),
                   .rst_in(sys_rst_pixel),

                   .write_valid_in(write_valid_in),
                   .write_addr_in(write_addr_in),
                   .write_object_in(write_object_in),
                   .write_valid_out(write_valid_out),

                   .read_valid_in(read_valid_in),
                   .read_addrs_in(read_addrs_in),
                   .read_objects_out(read_objects_out),
                   .read_valid_out(read_valid_out)
                 );

  // physics engine definition
  logic frame_start_in;
  enum logic [2:0] {IDLE, LOADING, COLLISION, UPDATING, SAVING} state_out;
  logic frame_end_out;

  logic load_signal_out;
  logic [`OBJ_ADDR_WIDTH-1:0] load_object_index_out [3:0];
  logic [`OBJ_WIDTH-1:0] load_object_data_in [3:0];

  logic save_signal_out;
  logic [`OBJ_ADDR_WIDTH-1:0] save_object_index_out;
  logic [`OBJ_WIDTH-1:0] save_object_data_out;

  physics_engine engine
                 (
                   .sys_clk(clk_pixel),
                   .sys_rst(sys_rst_pixel),
                   .frame_start_in(frame_start_in),
                   .state_out(state_out),
                   .frame_end_out(frame_end_out),

                   .load_signal_out(load_signal_out),
                   .load_object_index_out(load_object_index_out),
                   .load_object_data_in(load_object_data_in),

                   .save_signal_out(save_signal_out),
                   .save_object_index_out(save_object_index_out),
                   .save_object_data_out(save_object_data_out)
                 );


  logic is_obj_first_half;
  // BRAM integration
  always_ff @(posedge clk_pixel) // ff for buffering
  begin

    if(sys_rst_pixel) is_obj_first_half <= 0;
    else is_obj_first_half <= !is_obj_first_half;

    if (simul_mode)
    begin // IO from phys_engine
      write_valid_in <= save_signal_out | create_random_obj;
      if (save_signal_out)
      begin
        write_addr_in <= save_object_index_out;
        write_object_in <= save_object_data_out;
      end
      else if (create_random_obj)
      begin
        write_addr_in <= rd_idx;
        write_object_in <= random_obj;
      end
    end
    else
    begin // IO from draw & render
      write_valid_in <= 1'b0;
      // read_valid_in <= 1'b0;
    end

    if(is_memory_stable) begin
      // render reads
      if(is_obj_first_half) begin
        read_addrs_in <= {8'b0, 8'b1, 8'b10, 8'b11};
      end
      else begin
        read_addrs_in <= {8'b100, 8'b101, 8'b110, 8'b111};
      end
      
    end
    else begin
      // physics
      read_valid_in <= load_signal_out;
      if (load_signal_out)
      begin
        read_addrs_in[0] <= load_object_index_out[0];
        read_addrs_in[1] <= load_object_index_out[1];
        read_addrs_in[2] <= load_object_index_out[2];
        read_addrs_in[3] <= load_object_index_out[3];
      end
      if (read_valid_out)
      begin
        load_object_data_in[0] <= read_objects_out[0];
        load_object_data_in[1] <= read_objects_out[1];
        load_object_data_in[2] <= read_objects_out[2];
        load_object_data_in[3] <= read_objects_out[3];
      end
    end
  end

  // physics_engine integration
  assign frame_start_in = simul_mode && nf_hdmi && (!sw[14] || frame_count_hdmi[3:0] == 0); // slower framerate

  logic is_memory_stable;
  assign is_memory_stable = !simul_mode || (state_out == IDLE);
  assign led[15] = is_memory_stable;
  assign led[14] = simul_mode;
  assign led[13] = create_random_obj;


  // debugging obj0, obj1 ypos
  logic [15:0] obj0_pos_y, obj0_vel_y;
  logic [3:0] phys_ss0_an, phys_ss1_an;
  logic [6:0] phys_ss_c;

  seven_segment_controller phys_ssc(.clk_in(clk_pixel),
                                    .rst_in(sys_rst_pixel),
                                    .val_in({obj0_pos_y, obj0_vel_y}),
                                    .cat_out(phys_ss_c),
                                    .an_out({phys_ss0_an, phys_ss1_an}));


  logic frame_toggle;
  always_ff @(posedge clk_pixel)
  begin
    if(sys_rst_pixel)
    begin
      frame_toggle <= 1'b0;
    end
    else
      if(frame_start_in)
      begin
        frame_toggle <= ~frame_toggle;
      end
  end
  assign led[12] = frame_toggle;


  always_ff @(posedge clk_pixel)
  begin
    if(write_valid_in && write_addr_in == 0)
    begin
      obj0_pos_y <= write_object_in[47:32];
      obj0_vel_y <= write_object_in[15:0];
    end
  end

  // logic [15:0] prev_pos_y, prev_vel_y;
  // always_ff @(posedge clk_pixel)
  // begin
  //   if (sys_rst_pixel)
  //   begin
  //     prev_pos_y <= 0;
  //     prev_vel_y <= 0;
  //   end
  //   else
  //   begin
  //     if (create_random_obj)
  //     begin
  //       prev_pos_y <= pos_y;
  //       prev_vel_y <= vel_y;
  //     end
  //   end
  // end


  // debugging random objects
  logic create_random_obj;
  assign create_random_obj = btn[3];

  logic [15:0] rd_pos_xs[`OBJ_COUNT:0], rd_pos_ys[`OBJ_COUNT:0], rd_vel_xs[`OBJ_COUNT:0], rd_vel_ys[`OBJ_COUNT:0], rd_rads[`OBJ_COUNT:0];
  logic rd_is_static[`OBJ_COUNT:0];
  logic [`OBJ_WIDTH-1:0] random_obj;

  logic [2:0] rd_idx;
  logic [15:0] sd1, sd2;
  localparam RNG_A = 7603, RNG_C = 1557, RNG_MASK = 16'hFFFF;
  assign sd1 = (RNG_A * hcount_hdmi) & RNG_MASK + RNG_C;
  assign sd2 = (RNG_A * (vcount_hdmi ^ hcount_hdmi[3:0])) & RNG_MASK + RNG_C;

  always_ff @(posedge clk_pixel)
  begin
    if(create_random_obj)
    begin
      rd_pos_xs[rd_idx] <= {4'b0, sd1[11:0]};
      rd_pos_ys[rd_idx] <= {4'b0, ((RNG_A * sd1 + RNG_C) & RNG_MASK)};
      rd_vel_xs[rd_idx] <= {sd2[0], 5'b0, sd2[10:1]};
      rd_vel_ys[rd_idx] <= {sd2[13], 8'b0, sd2[15:11]};
      rd_rads[rd_idx] <= (sd1[7:0] ^ sd2[7:0]) & 16'h3FF + 16'h080;
      rd_is_static[rd_idx] <= (sd1[3] == 1'b1 && sd2[3] == 1'b1);

      random_obj <= 115'h1_000000000000_0000_0000_0000_0000 ^ (rd_is_static[rd_idx] << 112) ^ (rd_rads[rd_idx] << 64) ^ (rd_pos_xs[rd_idx] << 48) ^ (rd_pos_ys[rd_idx] << 32) ^ (rd_vel_xs[rd_idx] << 16) ^ rd_vel_ys[rd_idx];

      rd_idx <= rd_idx + 1;
    end
  end
  

  // logic [15:0] pos_y, vel_y; // both random
  // logic [`OBJ_WIDTH-1:0] random_obj;
  // assign pos_y = hcount_hdmi << 2;
  // assign vel_y = ~((hcount_hdmi[3:0] << 5) + (vcount_hdmi >> 3));
  // always_ff @(posedge clk_pixel)
  // begin
  //   if(create_random_obj)
  //   begin
  //     random_obj <= 115'h1_000000000a00_1900_0000_00a0_0000 + (pos_y << 32) + vel_y;
  //   end
  // end



  // object coordinate setting logic
  logic [86:0] obj_coord;
  always_comb
  begin
    if (btn[2])
    begin
      case (sw[7:6])
        2'b00:
          obj_coord = 87'b0;
        2'b01:
          obj_coord = {sw[2], sw[7:6], circle_coord};
        2'b10:
          obj_coord = {sw[2], sw[7:6], line_coord};
        2'b11:
          obj_coord = {sw[2], sw[7:6], rect_coord};
        default:
          obj_coord = 87'b0;
      endcase
    end
  end


  // HDMI video signal generator
  video_sig_gen vsg
                (
                  .pixel_clk_in(clk_pixel),
                  .rst_in(sys_rst_pixel),
                  .hcount_out(hcount_hdmi),
                  .vcount_out(vcount_hdmi),
                  .vs_out(vsync_hdmi),
                  .hs_out(hsync_hdmi),
                  .nf_out(nf_hdmi),
                  .ad_out(active_draw_hdmi),
                  .fc_out(frame_count_hdmi)
                );

    // input wire clk_in,
    // input wire valid_in,
    // input wire rst_in,
    // // parameters for up to four objects at a time being passed in from object storage
    // input wire [3:0] is_static,
    // // input wire [3:0][6:0] current_addresses,
    // input wire [3:0][1:0] id_bits,
    // input wire [3:0][47:0] params,
    // input wire [3:0][15:0] pos_x,
    // input wire [3:0][15:0] pos_y,

    // // pixel coordinate that we are querying
    // input wire [10:0] hcount_in,
    // input wire [9:0] vcount_in,

    // // resulting color
    // output logic [1:0] color_bits,

    // // write location to frame buffer
    // output logic [18:0] write_address,

    // // output logic busy_out, // todo remove
    // output logic valid_out

  logic [3:0] render_input_is_static;
  logic [3:0][1:0] render_input_id_bits;
  logic [3:0][47:0] render_input_params;
  logic [3:0][15:0] render_input_pos_x;
  logic [3:0][15:0] render_input_pos_y;
  logic [1:0] render_output_color_bits;
  logic [18:0] render_output_write_address;
  logic render_output_valid_out;

genvar render_index;
generate
  for(render_index = 0; render_index <= 3; render_index = render_index + 1) begin
    assign {render_input_is_static[render_index], 
            render_input_id_bits[render_index], 
            render_input_pos_x[render_index], 
            render_input_pos_y[render_index], 
            render_input_params[render_index]} 
            = read_objects_out[render_index];
  end
endgenerate

  logic dbg_valid_in;
  // logic [15:0] dbg_pos_x [3:0];
  // logic [15:0] dbg_pos_y [3:0];
  logic [47:0] dbg_params [3:0];
  logic [1:0] dbg_id_bits [3:0];

  logic dbg_is_shape_ready [3:0];
  logic dbg_is_shape_drawn [3:0];
  logic [10:0] dbg_x_in_1s [3:0];
  logic [10:0] dbg_x_in_2s [3:0];
  logic [9:0] dbg_y_in_1s [3:0];
  logic [9:0] dbg_y_in_2s [3:0];
  logic [83:0] dbg_obj_coord [3:0];
  logic dbg_in_shape_bits [3:0];

  assign dbg_valid_in = nf_hdmi;

  genvar dbg_i;
  generate 
    for(dbg_i=0; dbg_i<4; dbg_i=dbg_i+1) begin
      circle_converter dbg_ball_converter (
          .is_valid_in(dbg_id_bits[dbg_i] == 2'b01 && dbg_valid_in),
          .pos_x(rd_pos_xs[dbg_i]),
          .pos_y(rd_pos_ys[dbg_i]),
          .params({32'b0, rd_rads[dbg_i]}),
          .x_in_1(dbg_x_in_1s[dbg_i]),
          .y_in_1(dbg_y_in_1s[dbg_i]),
          .x_in_2(dbg_x_in_2s[dbg_i]),
          .y_in_2(dbg_y_in_2s[dbg_i]),
          .is_valid_out(dbg_is_shape_ready[dbg_i])
        );

      draw_circle dbg_ball(
        .valid_in(dbg_is_shape_ready[dbg_i]),
        .clk_in(clk_pixel),
        .rst_in(sys_rst_pixel),
        .hcount_in(hcount_hdmi),
        .vcount_in(vcount_hdmi),
        .x_in_1(dbg_x_in_1s[dbg_i]),
        .y_in_1(dbg_y_in_1s[dbg_i]),
        .x_in_2(dbg_x_in_2s[dbg_i]),
        .y_in_2(dbg_y_in_2s[dbg_i]),
        .circle_coord(dbg_obj_coord[dbg_i]),
        .in_circle(dbg_in_shape_bits[dbg_i]),
        .valid_out(dbg_is_shape_drawn[dbg_i])
      );
    end
  endgenerate

  logic [1:0] dbg_merged_bits, dbg_color_bits;
  assign dbg_merged_bits = dbg_in_shape_bits[0] | dbg_in_shape_bits[1] | dbg_in_shape_bits[2] | dbg_in_shape_bits[3];
  assign dbg_color_bits = (dbg_merged_bits == 2'b11) ? 2'b01 : dbg_merged_bits;


  // render render_objects
  // (
  //   .clk_in(clk_pixel),
  //   .valid_in(active_draw_hdmi && is_memory_stable && !vcount_hdmi[0]),
  //   .rst_in(sys_rst_pixel),
  //   .is_static(render_input_is_static),
  //   .id_bits(render_input_id_bits),
  //   .pos_x(render_input_pos_x),
  //   .pos_y(render_input_pos_y),
  //   .params(render_input_params),
  //   .hcount_in(hcount_hdmi),
  //   .vcount_in(vcount_hdmi),
  //   .color_bits(render_output_color_bits),
  //   .write_address(render_output_write_address),
  //   .valid_out(render_output_valid_out)
  // );

    logic [1:0] frame_buff_output;
    // port a for writing from render
    // port b for reading to hdmi
    xilinx_true_dual_port_read_first_2_clock_ram #(
    .RAM_WIDTH(2),                       // Specify RAM data width
    .RAM_DEPTH(640*480),                     // Specify RAM depth (number of entries)
    .RAM_PERFORMANCE("HIGH_PERFORMANCE"), // Select "HIGH_PERFORMANCE" or "LOW_LATENCY"
    .INIT_FILE("")                        // Specify name/location of RAM initialization file if using one (leave blank if not)
    ) render_frame_buffer (
    .addra(render_output_write_address),   // Port A address bus, width determined from RAM_DEPTH
    .addrb((hcount_hdmi >> 1) + 640 * (vcount_hdmi >> 1)),   // Port B address bus, width determined from RAM_DEPTH
    .dina(render_output_color_bits),     // Port A RAM input data, width determined from RAM_WIDTH
    .dinb(),     // Port B RAM input data, width determined from RAM_WIDTH
    .clka(clk_pixel),     // Port A clock
    .clkb(clk_pixel),     // Port B clock
    .wea(render_output_valid_out),       // Port A write enable
    .web(0),       // Port B write enable
    .ena(1),       // Port A RAM Enable, for additional power savings, disable port when not in use
    .enb(1),       // Port B RAM Enable, for additional power savings, disable port when not in use
    .rsta(sys_rst_pixel),     // Port A output reset (does not affect memory contents)
    .rstb(sys_rst_pixel),     // Port B output reset (does not affect memory contents)
    .regcea(1), // Port A output register enable
    .regceb(), // Port B output register enable
    .douta(),   // Port A RAM output data, width determined from RAM_WIDTH
    .doutb(frame_buff_output)    // Port B RAM output data, width determined from RAM_WIDTH
  );


  // Video Mux: select from the different display modes based on switch values
  //used with switches for display selections
  logic [1:0] display_choice;
  logic [1:0] target_choice;

  assign display_choice = sw[5:4];
  assign target_choice =  sw[7:6];

  //choose what to display from the camera:
  // * 'b00:  normal camera out
  // * 'b01:  selected channel image in grayscale
  // * 'b10:  masked pixel (all on if 1, all off if 0)
  // * 'b11:  chroma channel with mask overtop as magenta
  //
  //then choose what to use with center of mass:
  // * 'b00: nothing
  // * 'b01: crosshair
  // * 'b10: sprite on top
  // * 'b11: nothing

  logic [7:0] fb_red_delayed_ps2;
  pipeline #(
             .WIDTH(8), .STAGES(4))
           fb_red_pipeline_ps2(
             .clk_pixel(clk_pixel),
             .signal(fb_red),
             //.stages(4),
             .delayed_signal(fb_red_delayed_ps2)
           );

  logic [7:0] fb_green_delayed_ps2;
  pipeline #(
             .WIDTH(8), .STAGES(4))
           fb_green_pipeline_ps2(
             .clk_pixel(clk_pixel),
             .signal(fb_green),
             //.stages(4),
             .delayed_signal(fb_green_delayed_ps2)
           );

  logic [7:0] fb_blue_delayed_ps2;
  pipeline #(
             .WIDTH(8), .STAGES(4))
           fb_blue_pipeline_ps2(
             .clk_pixel(clk_pixel),
             .signal(fb_blue),
             //.stages(4),
             .delayed_signal(fb_blue_delayed_ps2)
           );

  logic [7:0] y_delayed_ps6;
  pipeline #(
             .WIDTH(8), .STAGES(1))
           y_pipeline_ps6(
             .clk_pixel(clk_pixel),
             .signal(y),
             //.stages(1),
             .delayed_signal(y_delayed_ps6)
           );

  logic [7:0] selected_channel_delayed_ps5;
  pipeline #(
             .WIDTH(8), .STAGES(1))
           selected_channel_pipeline_ps5(
             .clk_pixel(clk_pixel),
             .signal(selected_channel),
             //.stages(1),
             .delayed_signal(selected_channel_delayed_ps5)
           );


/*
module video_mux (
  // input wire [1:0] bg_in, //regular video
  input wire [1:0] target_in, //regular video
  // input wire [23:0] camera_pixel_in, //16 bits from camera 5:6:5
  // input wire [7:0] camera_y_in,  //y channel of ycrcb camera conversion
  // input wire [7:0] channel_in, //the channel from selection module
  // input wire thresholded_pixel_in, //
  input wire [1:0] frame_buff_out,
  input wire rect_pixel_in,
  input wire circle_pixel_in,
  input wire line_pixel_in,
  output logic [23:0] pixel_out
);
*/
  video_mux mvm(
              // .bg_in(display_choice), //choose background
              .target_in(target_choice), //choose target
              // .camera_pixel_in({fb_red_delayed_ps2, fb_green_delayed_ps2, fb_blue_delayed_ps2}), //TODO: needs (PS2)
              // .camera_y_in(y_delayed_ps6), //luminance TODO: needs (PS6)
              // .channel_in(selected_channel_delayed_ps5), //current channel being drawn TODO: needs (PS5)
              // .thresholded_pixel_in(mask), //one bit mask signal TODO: needs (PS4)
              .frame_buff_out(dbg_color_bits), //output from frame buffer
              .rect_pixel_in(in_rect), //TODO: needs (PS9) maybe?
              .circle_pixel_in(in_circle),
              .line_pixel_in(in_line),
              .pixel_out({red,green,blue}) //output to tmds
            );

  // HDMI Output: just like before!

  logic [9:0] tmds_10b [0:2]; //output of each TMDS encoder!
  logic       tmds_signal [2:0]; //output of each TMDS serializer!

  //three tmds_encoders (blue, green, red)
  //note green should have no control signal like red
  //the blue channel DOES carry the two sync signals:
  //  * control_in[0] = horizontal sync signal
  //  * control_in[1] = vertical sync signal

  tmds_encoder tmds_red(
                 .clk_in(clk_pixel),
                 .rst_in(sys_rst_pixel),
                 .data_in(red),
                 .control_in(2'b0),
                 .ve_in(active_draw_hdmi),
                 .tmds_out(tmds_10b[2]));

  tmds_encoder tmds_green(
                 .clk_in(clk_pixel),
                 .rst_in(sys_rst_pixel),
                 .data_in(green),
                 .control_in(2'b0),
                 .ve_in(active_draw_hdmi),
                 .tmds_out(tmds_10b[1]));

  tmds_encoder tmds_blue(
                 .clk_in(clk_pixel),
                 .rst_in(sys_rst_pixel),
                 .data_in(blue),
                 .control_in({vsync_hdmi,hsync_hdmi}),
                 .ve_in(active_draw_hdmi),
                 .tmds_out(tmds_10b[0]));


  //three tmds_serializers (blue, green, red):
  //MISSING: two more serializers for the green and blue tmds signals.
  tmds_serializer red_ser(
                    .clk_pixel_in(clk_pixel),
                    .clk_5x_in(clk_5x),
                    .rst_in(sys_rst_pixel),
                    .tmds_in(tmds_10b[2]),
                    .tmds_out(tmds_signal[2]));
  tmds_serializer green_ser(
                    .clk_pixel_in(clk_pixel),
                    .clk_5x_in(clk_5x),
                    .rst_in(sys_rst_pixel),
                    .tmds_in(tmds_10b[1]),
                    .tmds_out(tmds_signal[1]));
  tmds_serializer blue_ser(
                    .clk_pixel_in(clk_pixel),
                    .clk_5x_in(clk_5x),
                    .rst_in(sys_rst_pixel),
                    .tmds_in(tmds_10b[0]),
                    .tmds_out(tmds_signal[0]));

  //output buffers generating differential signals:
  //three for the r,g,b signals and one that is at the pixel clock rate
  //the HDMI receivers use recover logic coupled with the control signals asserted
  //during blanking and sync periods to synchronize their faster bit clocks off
  //of the slower pixel clock (so they can recover a clock of about 742.5 MHz from
  //the slower 74.25 MHz clock)
  OBUFDS OBUFDS_blue (.I(tmds_signal[0]), .O(hdmi_tx_p[0]), .OB(hdmi_tx_n[0]));
  OBUFDS OBUFDS_green(.I(tmds_signal[1]), .O(hdmi_tx_p[1]), .OB(hdmi_tx_n[1]));
  OBUFDS OBUFDS_red  (.I(tmds_signal[2]), .O(hdmi_tx_p[2]), .OB(hdmi_tx_n[2]));
  OBUFDS OBUFDS_clock(.I(clk_pixel), .O(hdmi_clk_p), .OB(hdmi_clk_n));


  // Nothing To Touch Down Here:
  // register writes to the camera

  // The OV5640 has an I2C bus connected to the board, which is used
  // for setting all the hardware settings (gain, white balance,
  // compression, image quality, etc) needed to start the camera up.
  // We've taken care of setting these all these values for you:
  // "rom.mem" holds a sequence of bytes to be sent over I2C to get
  // the camera up and running, and we've written a design that sends
  // them just after a reset completes.

  // If the camera is not giving data, press your reset button.

  logic  busy, bus_active;
  logic  cr_init_valid, cr_init_ready;

  logic  recent_reset;
  always_ff @(posedge clk_camera)
  begin
    if (sys_rst_camera)
    begin
      recent_reset <= 1'b1;
      cr_init_valid <= 1'b0;
    end
    else if (recent_reset)
    begin
      cr_init_valid <= 1'b1;
      recent_reset <= 1'b0;
    end
    else if (cr_init_valid && cr_init_ready)
    begin
      cr_init_valid <= 1'b0;
    end
  end

  logic [23:0] bram_dout;
  logic [7:0]  bram_addr;

  // ROM holding pre-built camera settings to send
  xilinx_single_port_ram_read_first
    #(
      .RAM_WIDTH(24),
      .RAM_DEPTH(256),
      .RAM_PERFORMANCE("HIGH_PERFORMANCE"),
      .INIT_FILE("rom.mem")
    ) registers
    (
      .addra(bram_addr),     // Address bus, width determined from RAM_DEPTH
      .dina(24'b0),          // RAM input data, width determined from RAM_WIDTH
      .clka(clk_camera),     // Clock
      .wea(1'b0),            // Write enable
      .ena(1'b1),            // RAM Enable, for additional power savings, disable port when not in use
      .rsta(sys_rst_camera), // Output reset (does not affect memory contents)
      .regcea(1'b1),         // Output register enable
      .douta(bram_dout)      // RAM output data, width determined from RAM_WIDTH
    );

  logic [23:0] registers_dout;
  logic [7:0]  registers_addr;
  assign registers_dout = bram_dout;
  assign bram_addr = registers_addr;

  logic       con_scl_i, con_scl_o, con_scl_t;
  logic       con_sda_i, con_sda_o, con_sda_t;

  // NOTE these also have pullup specified in the xdc file!
  // access our inouts properly as tri-state pins
  IOBUF IOBUF_scl (.I(con_scl_o), .IO(i2c_scl), .O(con_scl_i), .T(con_scl_t) );
  IOBUF IOBUF_sda (.I(con_sda_o), .IO(i2c_sda), .O(con_sda_i), .T(con_sda_t) );

  // provided module to send data BRAM -> I2C
  camera_registers crw
                   (.clk_in(clk_camera),
                    .rst_in(sys_rst_camera),
                    .init_valid(cr_init_valid),
                    .init_ready(cr_init_ready),
                    .scl_i(con_scl_i),
                    .scl_o(con_scl_o),
                    .scl_t(con_scl_t),
                    .sda_i(con_sda_i),
                    .sda_o(con_sda_o),
                    .sda_t(con_sda_t),
                    .bram_dout(registers_dout),
                    .bram_addr(registers_addr));

  // a handful of debug signals for writing to registers
  assign led[0] = crw.bus_active;
  assign led[1] = cr_init_valid;
  assign led[2] = cr_init_ready;
  // assign led[15:3] = 0;

endmodule // top_level


`default_nettype wire
