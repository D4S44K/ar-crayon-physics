module render
  (
    input wire clk_in,
    input wire valid_in,
    input wire rst_in,
    // parameters for up to four objects at a time being passed in from object storage
    input wire [3:0] is_static,
    // input wire [3:0][6:0] current_addresses,
    input wire [3:0][1:0] id_bits,
    input wire [3:0][47:0] params,
    input wire [3:0][15:0] pos_x,
    input wire [3:0][15:0] pos_y,

    // pixel coordinate that we are querying
    input wire [10:0] hcount_in,
    input wire [9:0] vcount_in,

    // resulting color
    output logic [1:0] color_bits,

    // write location to frame buffer
    output logic [18:0] write_address,

    // output logic busy_out, // todo remove
    output logic valid_out
  );

  localparam STATIC_COLOR = 24'h11_11_11;
  localparam NOT_STATIC_COLOR = 24'h77_77_77;

  logic [11:0][10:0] x_in_1s;
  logic [11:0][9:0] y_in_1s;
  logic [11:0][10:0] x_in_2s;
  logic [11:0][9:0] y_in_2s;
  // 00: black, 01: color it static, 10: color it movable, 11: n/a right now
  logic [3:0][23:0] colors;
  logic [11:0] in_shape_bits;
  logic [11:0][83:0] obj_coord;
  logic [11:0] is_shape_ready;
  logic [11:0] is_shape_drawn;

  genvar i;
  generate
    begin
      for(i=0; i<4; i++)
      begin
        draw_circle  ball(
                       .valid_in(is_shape_ready[i]),
                       .clk_in(clk_in),
                       .rst_in(rst_in),
                       .hcount_in(hcount_in),
                       .vcount_in(vcount_in),
                       .x_in_1(x_in_1s[i]),
                       .y_in_1(y_in_1s[i]),
                       .x_in_2(x_in_2s[i]),
                       .y_in_2(y_in_2s[i]),
                       .circle_coord(obj_coord[i]),
                       .in_circle(in_shape_bits[i]),
                       .valid_out(is_shape_drawn[i])
                     );

        circle_converter ball_converter (
                           // .is_static(is_static[0]),
                           .is_valid_in(id_bits[i] == 2'b01 && valid_in),
                           .pos_x(pos_x[i]),
                           .pos_y(pos_y[i]),
                           .params(params[i]),
                           .x_in_1(x_in_1s[i]),
                           .y_in_1(y_in_1s[i]),
                           .x_in_2(x_in_2s[i]),
                           .y_in_2(y_in_2s[i]),
                           .is_valid_out(is_shape_ready[i])
                         );
      end
    end
  endgenerate

  generate
    for(i=0; i<4; i++)
    begin
      draw_line  line(
                   .valid_in(is_shape_ready[4+i] ),
                   .clk_in(clk_in),
                   .rst_in(rst_in),
                   .hcount_in(hcount_in),
                   .vcount_in(vcount_in),
                   .x_in_1(x_in_1s[4+i]),
                   .y_in_1(y_in_1s[4+i]),
                   .x_in_2(x_in_2s[4+i]),
                   .y_in_2(y_in_2s[4+i]),
                   .line_coord(obj_coord[4+i]),
                   .in_line(in_shape_bits[4+i]),
                   .valid_out(is_shape_drawn[4+i])
                 );

      line_converter line_converter (
                       // .is_static(is_static[0]),
                       .is_valid_in(id_bits[i] == 2'b10 && valid_in),
                       .pos_x(pos_x[i]),
                       .pos_y(pos_y[i]),
                       .params(params[i]),
                       .x_in_1(x_in_1s[4+i]),
                       .y_in_1(y_in_1s[4+i]),
                       .x_in_2(x_in_2s[4+i]),
                       .y_in_2(y_in_2s[4+i]),
                       .is_valid_out(is_shape_ready[4+i])
                     );
    end
  endgenerate

  generate
    for(i=0; i<4; i++)
    begin
      draw_rectangle  rect(
                        .valid_in(is_shape_ready[8+i]),
                        .clk_in(clk_in),
                        .rst_in(rst_in),
                        .hcount_in(hcount_in),
                        .vcount_in(vcount_in),
                        .x_in_1(x_in_1s[8+i]),
                        .y_in_1(y_in_1s[8+i]),
                        .x_in_2(x_in_2s[8+i]),
                        .y_in_2(y_in_2s[8+i]),
                        .rect_coord(obj_coord[8+i]),
                        .in_rect(in_shape_bits[8+i]),
                        .valid_out(is_shape_drawn[8+i])
                      );

      rect_converter rect_converter (
                       // .is_static(is_static[0]),
                       .is_valid_in(id_bits[i] ==2'b11 && valid_in),
                       .pos_x(pos_x[i]),
                       .pos_y(pos_y[i]),
                       .params(params[i]),
                       .x_in_1(x_in_1s[8+i]),
                       .y_in_1(y_in_1s[8+i]),
                       .x_in_2(x_in_2s[8+i]),
                       .y_in_2(y_in_2s[8+i]),
                       .is_valid_out(is_shape_ready[8+i])
                     );
    end
  endgenerate


  logic [3:0] held_in_shape_bits;
  logic [4:0][18:0] held_write_address;
  logic [18:0] cycle_delay_write_address;
  // logic [4:0][3:0] held_valid;
  logic [5:0][3:0][1:0] held_id_bits_set_1;
  logic [4:0][3:0][1:0] held_id_bits_set_2;
  logic [5:0][3:0] held_static_bits_set_1;
  logic [4:0][3:0] held_static_bits_set_2;
  logic [4:0] held_is_second_set;
  logic [3:0] current_in_shape_bits;
  logic [1:0] final_color_bit;
  logic is_second_set;

  // determines whether the pointeger is in the second set of shapes
  always_comb
  begin
    for(integer obj_num = 0; obj_num < 4; obj_num = obj_num + 1)
    begin
      case(held_id_bits_set_2[obj_num])
        2'b00:
          current_in_shape_bits[obj_num] = 0;
        2'b01:
          current_in_shape_bits[obj_num] = in_shape_bits[obj_num];
        2'b10:
          current_in_shape_bits[obj_num] = in_shape_bits[obj_num + 4];
        2'b11:
          current_in_shape_bits[obj_num] = in_shape_bits[obj_num+8];
        default:
          current_in_shape_bits[obj_num] = 0;
      endcase
    end
  end

  always_ff@(posedge clk_in)
  begin
    if(rst_in)
    begin
      valid_out <= 0;
      held_in_shape_bits <= 0;
      is_second_set <= 0;
      held_is_second_set <= 0;
      held_id_bits_set_1 <= 0;
      held_id_bits_set_2 <= 0;
      held_static_bits_set_1 <= 0;
      held_static_bits_set_2 <= 0;
      color_bits <= 0;
      cycle_delay_write_address <= 0;
      held_write_address <= 0;
    end
    else if(valid_in)
    begin
      is_second_set <= !is_second_set;
      for(integer i = 0; i <= 3; i = i + 1)
      begin
        held_is_second_set[i + 1] <= held_is_second_set[i];
        held_id_bits_set_1[i + 1] <= held_id_bits_set_1[i];
        held_id_bits_set_2[i + 1] <= held_id_bits_set_2[i];
        held_write_address[i + 1] <= held_write_address[i];
        held_static_bits_set_1[i + 1] <= held_static_bits_set_1[i];
        held_static_bits_set_2[i + 1] <= held_static_bits_set_2[i];
      end
      held_is_second_set[0] <= is_second_set;
      if(!is_second_set)
        held_id_bits_set_1[0] <= id_bits;
      else
        held_id_bits_set_2[0] <= id_bits;
      if(is_second_set)
        held_static_bits_set_2[0] <= is_static;
      else
        held_static_bits_set_1[0] <= is_static;
      held_static_bits_set_1[5] <= held_static_bits_set_1[4];
      held_id_bits_set_1[5] <= held_id_bits_set_1[4];
      held_write_address[0] <= (hcount_in >> 1) + (640 * (vcount_in >> 1));

      if(!held_is_second_set[4])
      begin
        cycle_delay_write_address <= held_write_address[4];
        for(integer obj_num = 0; obj_num < 4; obj_num = obj_num + 1)
        begin
          case(held_id_bits_set_1[5][obj_num])
            2'b00:
              held_in_shape_bits[obj_num] <= 0;
            2'b01:
              held_in_shape_bits[obj_num] <= in_shape_bits[obj_num];
            2'b10:
              held_in_shape_bits[obj_num] <= in_shape_bits[obj_num + 4];
            2'b11:
              held_in_shape_bits[obj_num] <= in_shape_bits[obj_num+8];
            default:
              held_in_shape_bits[obj_num] <= 0;
          endcase
        end
        valid_out <= 0;

      end
      else
      begin
        if(held_in_shape_bits[0])
          color_bits <= held_static_bits_set_1[0] ? 2'b10 : 2'b01;
        else if(held_in_shape_bits[1])
          color_bits <= held_static_bits_set_1[1] ? 2'b10 : 2'b01;
        else if(held_in_shape_bits[2])
          color_bits <= held_static_bits_set_1[2] ? 2'b10 : 2'b01;
        else if(held_in_shape_bits[3])
          color_bits <= held_static_bits_set_1[3] ? 2'b10 : 2'b01;
        else if(current_in_shape_bits[0])
          color_bits <= held_static_bits_set_2[0] ? 2'b10 : 2'b01;
        else if(current_in_shape_bits[1])
          color_bits <= held_static_bits_set_2[1] ? 2'b10 : 2'b01;
        else if(current_in_shape_bits[2])
          color_bits <= held_static_bits_set_2[2] ? 2'b10 : 2'b01;
        else if(current_in_shape_bits[3])
          color_bits <= held_static_bits_set_2[3] ? 2'b10 : 2'b01;
        else
          color_bits <= 2'b11;
        valid_out <= 1;
        write_address <= cycle_delay_write_address;

      end

    end
  end
endmodule
