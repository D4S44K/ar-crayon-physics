// `default_nettype none
// module update_collision_vel #(OBJ_WIDTH=128, PART_WIDTH=66, DF=32, SF=16)(
//     input wire sys_clk,
//     input wire sys_rst,
//     input wire data_valid_in,
//     input wire [OBJ_WIDTH-1:0] obj_a,
//     input wire [OBJ_WIDTH-1:0] obj_b,
//     input wire [2:0] a_part_index,
//     input wire [2:0] b_part_index

//     output wire data_valid_out,
//     output wire [SF-1:0] obj_a_rv_x,
//     output wire [SF-1:0] obj_a_rv_y,
//     output wire [SF-1:0] obj_b_rv_x,
//     output wire [SF-1:0] obj_b_rv_y
//   );
//   // should be completed in 16 cycles


// endmodule
