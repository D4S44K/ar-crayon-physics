module video_sig_gen
  #(
     parameter ACTIVE_H_PIXELS = 1280,
     parameter H_FRONT_PORCH = 110,
     parameter H_SYNC_WIDTH = 40,
     parameter H_BACK_PORCH = 220,
     parameter ACTIVE_LINES = 720,
     parameter V_FRONT_PORCH = 5,
     parameter V_SYNC_WIDTH = 5,
     parameter V_BACK_PORCH = 20,
     parameter FPS = 60)
   (
     input wire pixel_clk_in,
     input wire rst_in,
     output logic [$clog2(TOTAL_PIXELS)-1:0] hcount_out,
     output logic [$clog2(TOTAL_LINES)-1:0] vcount_out,
     output logic vs_out, //vertical sync out
     output logic hs_out, //horizontal sync out
     output logic ad_out,
     output logic nf_out, //single cycle enable signal
     output logic [5:0] fc_out); //frame

  localparam TOTAL_PIXELS = ACTIVE_H_PIXELS + H_FRONT_PORCH + H_SYNC_WIDTH + H_BACK_PORCH;
  localparam TOTAL_LINES = ACTIVE_LINES + V_FRONT_PORCH + V_SYNC_WIDTH + V_BACK_PORCH;

  logic fresh_start;

  always_ff @(posedge pixel_clk_in)
  begin
    if (rst_in)
    begin
      // reset all output and state
      fresh_start <= 1;
      hcount_out <= 0;
      vcount_out <= 0;
      fc_out <= 0;
    end
    else
    begin
      if (fresh_start)
      begin
        fresh_start <= 0;
        hcount_out <= 0;
        vcount_out <= 0;
      end
      else
      begin
        if (hcount_out == TOTAL_PIXELS - 1)
        begin
          hcount_out <= 0;
          if (vcount_out == TOTAL_LINES - 1)
          begin
            vcount_out <= 0;
            if (fc_out == FPS - 1)
            begin
              fc_out <= 0;
            end
            else
            begin
              fc_out <= fc_out + 1;
            end
          end
          else
          begin
            vcount_out <= vcount_out + 1;
          end
        end
        else
        begin
          hcount_out <= hcount_out + 1;
          vcount_out <= vcount_out;
        end
      end
    end
  end

  always_comb
  begin
    if (rst_in)
    begin
      vs_out = 1'b0;
      hs_out = 1'b0;
      ad_out = 1'b0;
      nf_out = 1'b0;
    end
    else
    begin
      if (hcount_out < ACTIVE_H_PIXELS)
      begin
        if (vcount_out < ACTIVE_LINES)
        begin
          hs_out = 1'b0;
          ad_out = 1'b1;
        end
      end
      else if (hcount_out < ACTIVE_H_PIXELS + H_FRONT_PORCH)
      begin
        hs_out = 1'b0;
        ad_out = 1'b0;
      end
      else if (hcount_out < ACTIVE_H_PIXELS + H_FRONT_PORCH + H_SYNC_WIDTH)
      begin
        hs_out = 1'b1;
        ad_out = 1'b0;
      end
      else if (hcount_out < TOTAL_PIXELS)
      begin
        hs_out = 1'b0;
        ad_out = 1'b0;
      end
      else
      begin
        // should not happen
      end

      if (vcount_out < ACTIVE_LINES)
      begin
        vs_out = 1'b0;
      end
      else if (vcount_out < ACTIVE_LINES + V_FRONT_PORCH)
      begin
        vs_out = 1'b0;
      end
      else if (vcount_out < ACTIVE_LINES + V_FRONT_PORCH + V_SYNC_WIDTH)
      begin
        vs_out = 1'b1;
      end
      else if (vcount_out < TOTAL_LINES)
      begin
        vs_out = 1'b0;
      end
      else
      begin
        // should not happen
      end

      if (hcount_out == ACTIVE_H_PIXELS && vcount_out == ACTIVE_LINES)
      begin
        nf_out = 1'b1;
      end
      else
      begin
        nf_out = 1'b0;
      end
    end
  end

endmodule
