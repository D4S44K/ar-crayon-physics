`default_nettype none
module get_part_collision #(PART_WIDTH=66, DF=32, SF=16)(
    input wire sys_clk,
    input wire sys_rst,
    input wire data_valid_in,
    input wire [PART_WIDTH-1:0] part_a,
    input wire [PART_WIDTH-1:0] part_b,
    input wire [SF-1:0] rv_x,
    input wire [SF-1:0] rv_y,

    output wire data_valid_out,
    output wire [DF-1:0] col_time,
  );

  // should be completed in 50 cycles


endmodule
